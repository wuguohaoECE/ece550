module thirty_two_bit_or(out, A, B);

	parameter SIZE = 32;
	input [SIZE-1:0] A,B;
	
	
	output [SIZE-1:0] out;
	
	or or_0(out[0], A[0], B[0]);
	or or_1(out[1], A[1], B[1]);
	or or_2(out[2], A[2], B[2]);
	or or_3(out[3], A[3], B[3]);
	or or_4(out[4], A[4], B[4]);
	or or_5(out[5], A[5], B[5]);
	or or_6(out[6], A[6], B[6]);
	or or_7(out[7], A[7], B[7]);
	or or_8(out[8], A[8], B[8]);
	or or_9(out[9], A[9], B[9]);
	or or_10(out[10], A[10], B[10]);
	or or_11(out[11], A[11], B[11]);
	or or_12(out[12], A[12], B[12]);
	or or_13(out[13], A[13], B[13]);
	or or_14(out[14], A[14], B[14]);
	or or_15(out[15], A[15], B[15]);
	or or_16(out[16], A[16], B[16]);
	or or_17(out[17], A[17], B[17]);
	or or_18(out[18], A[18], B[18]);
	or or_19(out[19], A[19], B[19]);
	or or_20(out[20], A[20], B[20]);
	or or_21(out[21], A[21], B[21]);
	or or_22(out[22], A[22], B[22]);
	or or_23(out[23], A[23], B[23]);
	or or_24(out[24], A[24], B[24]);
	or or_25(out[25], A[25], B[25]);
	or or_26(out[26], A[26], B[26]);
	or or_27(out[27], A[27], B[27]);
	or or_28(out[28], A[28], B[28]);
	or or_29(out[29], A[29], B[29]);
	or or_30(out[30], A[30], B[30]);
	or or_31(out[31], A[31], B[31]);

endmodule