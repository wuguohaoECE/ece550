module thirty_two_bit_splitter(in, Out);

	parameter SIZE = 32;
	input in;
	
	
	output [SIZE-1:0] Out;
	assign Out[0] = in;
	assign Out[1] = in;
	assign Out[2] = in;
	assign Out[3] = in;
	assign Out[4] = in;
	assign Out[5] = in;
	assign Out[6] = in;
	assign Out[7] = in;
	assign Out[8] = in;
	assign Out[9] = in;
	assign Out[10] = in;
	assign Out[11] = in;
	assign Out[12] = in;
	assign Out[13] = in;
	assign Out[14] = in;
	assign Out[15] = in;
	assign Out[16] = in;
	assign Out[17] = in;
	assign Out[18] = in;
	assign Out[19] = in;
	assign Out[20] = in;
	assign Out[21] = in;
	assign Out[22] = in;
	assign Out[23] = in;
	assign Out[24] = in;
	assign Out[25] = in;
	assign Out[26] = in;
	assign Out[27] = in;
	assign Out[28] = in;
	assign Out[29] = in;
	assign Out[30] = in;
	assign Out[31] = in;

endmodule